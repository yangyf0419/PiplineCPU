// rom_test4.v
// test UART
//`timescale 1ns/1ps

module ROM_4 (addr,data);
    input [31:0] addr;
    output [31:0] data;
    reg [31:0] data;
    localparam ROM_SIZE = 32;
    reg [31:0] ROM_DATA[ROM_SIZE-1:0];

    always@(*)
        case(addr[17:2])   //Address Must Be Word Aligned.
            16'd0: data <= {6'b000010, 26'b00000000000000000000001100};
            16'd1: data <= {6'b000010, 26'b00000000000000000000010001};
            16'd2: data <= {6'b000010, 26'b00000000000000000000010010};
            16'd3: data <= {6'b101011, 5'b11001, 5'b10111, 16'b0000000000100000};
            16'd4: data <= {6'b100011, 5'b11001, 5'b01000, 16'b0000000000100000};
            16'd5: data <= {6'b001100, 5'b01000, 5'b01001, 16'b0000000000001000};
            16'd6: data <= {6'b000100, 5'b01001, 5'b00000, 16'b1111111111111101};
            16'd7: data <= {6'b001100, 5'b01000, 5'b01000, 16'b1111111111111100};
            16'd8: data <= {6'b101011, 5'b11001, 5'b01000, 16'b0000000000100000};
            16'd9: data <= {6'b100011, 5'b11001, 5'b00100, 16'b0000000000011100};
            16'd10: data <= {6'b101011, 5'b11001, 5'b00100, 16'b0000000000001100};
            16'd11: data <= {6'b000010, 26'b00000000000000000000000011};
            16'd12: data <= {6'b001000, 5'b00000, 5'b11111, 16'b0000000000001100};
            16'd13: data <= {6'b001111, 5'b00000, 5'b11011, 16'b1000000000000000};
            16'd14: data <= {6'b001111, 5'b00000, 5'b11001, 16'b0100000000000000};
            16'd15: data <= {6'b001000, 5'b00000, 5'b10111, 16'b0000000000000010};
            16'd16: data <= {6'b000000, 5'b11111, 5'b00000, 5'b00000, 5'b00000, 6'b001000};
            16'd17: data <= {6'b000000, 5'b11010, 5'b00000, 5'b00000, 5'b00000, 6'b001000};
            16'd18: data <= {6'b000000, 5'b11010, 5'b00000, 5'b00000, 5'b00000, 6'b001000};
            default: data <= 32'h80000000;
        endcase
endmodule


