// rom_test6.v
// test CPU
//`timescale 1ns/1ps

module ROM_6 (addr,data);
    input [31:0] addr;
    output [31:0] data;
    reg [31:0] data;
    localparam ROM_SIZE = 32;
    reg [31:0] ROM_DATA[ROM_SIZE-1:0];

    always@(*)
        case(addr[17:2])   //Address Must Be Word Aligned.
            16'd0: data <= {6'b000010, 26'b00000000000000000000011000};
            16'd1: data <= {6'b000010, 26'b00000000000000000000011011};
            16'd2: data <= {6'b000010, 26'b00000000000000000000011100};
            16'd3: data <= {6'b001000, 5'b00000, 5'b00100, 16'b0011000000111001};
            16'd4: data <= {6'b101011, 5'b11001, 5'b00100, 16'b0000000000001100};
            16'd5: data <= {6'b001001, 5'b00000, 5'b00101, 16'b1101010000110001};
            16'd6: data <= {6'b101011, 5'b11001, 5'b00101, 16'b0000000000001100};
            16'd7: data <= {6'b000000, 5'b00000, 5'b00101, 5'b00110, 5'b10000, 6'b000000};
            16'd8: data <= {6'b101011, 5'b11001, 5'b00110, 16'b0000000000001100};
            16'd9: data <= {6'b000000, 5'b00000, 5'b00110, 5'b00111, 5'b10000, 6'b000011};
            16'd10: data <= {6'b101011, 5'b11001, 5'b00111, 16'b0000000000001100};
            16'd11: data <= {6'b000100, 5'b00111, 5'b00101, 16'b0000000000000001};
            16'd12: data <= {6'b001111, 5'b00000, 5'b00100, 16'b1101010010011001};
            16'd13: data <= {6'b000000, 5'b00110, 5'b00100, 5'b01000, 5'b00000, 6'b100000};
            16'd14: data <= {6'b101011, 5'b11001, 5'b01000, 16'b0000000000001100};
            16'd15: data <= {6'b000000, 5'b00000, 5'b01000, 5'b01001, 5'b01000, 6'b000011};
            16'd16: data <= {6'b101011, 5'b11001, 5'b01001, 16'b0000000000001100};
            16'd17: data <= {6'b001000, 5'b00000, 5'b01010, 16'b1100111111000111};
            16'd18: data <= {6'b101011, 5'b11001, 5'b01010, 16'b0000000000001100};
            16'd19: data <= {6'b000000, 5'b00100, 5'b01010, 5'b00010, 5'b00000, 6'b101010};
            16'd20: data <= {6'b101011, 5'b11001, 5'b00010, 16'b0000000000001100};
            16'd21: data <= {6'b000000, 5'b00100, 5'b01010, 5'b00011, 5'b00000, 6'b101011};
            16'd22: data <= {6'b101011, 5'b11001, 5'b00011, 16'b0000000000001100};
            16'd23: data <= {6'b000010, 26'b00000000000000000000010111};
            16'd24: data <= {6'b001000, 5'b00000, 5'b11111, 16'b0000000000001100};
            16'd25: data <= {6'b001111, 5'b00000, 5'b11001, 16'b0100000000000000};
            16'd26: data <= {6'b000000, 5'b11111, 5'b00000, 5'b00000, 5'b00000, 6'b001000};
            16'd27: data <= {6'b000000, 5'b11010, 5'b00000, 5'b00000, 5'b00000, 6'b001000};
            16'd28: data <= {6'b000000, 5'b11010, 5'b00000, 5'b00000, 5'b00000, 6'b001000};
            
            default: data <= 32'h80000000;
        endcase
endmodule


