// hazard_units.v
// hazard_detection_unit, bypassing_unit


module hazard_detection_unit();