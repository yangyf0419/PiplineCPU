`timescale 1ns/1ns

//指令存储器

module ROM1 (addr,data);
input [31:0] addr;
output [31:0] data;
reg [31:0] data;

always@(*)
	case(addr[8:2])	//Address Must Be Word Aligned.
		7'd0: data <= {6'b001000, 5'b00000, 5'b10001, 16'b0000000000000001};
		7'd1: data <= {6'b001000, 5'b00000, 5'b10010, 16'b0000000000000010};
		7'd2: data <= {6'b001000, 5'b00000, 5'b10011, 16'b0000000000000011};
		7'd3: data <= {6'b100011, 5'b00000, 5'b10001, 16'b0000000000000000};
		7'd4: data <= {6'b100011, 5'b00000, 5'b10010, 16'b0000000000000100};
		7'd5: data <= {6'b100011, 5'b00000, 5'b10011, 16'b0000000000001000};
		7'd6: data <= {6'b000000, 5'b10001, 5'b10010, 5'b01000, 5'b00000, 6'b100000};
		7'd7: data <= {6'b000000, 5'b10001, 5'b10011, 5'b01001, 5'b00000, 6'b100000};
		7'd8: data <= {6'b000000, 5'b01000, 5'b01001, 5'b01000, 5'b00000, 6'b100000};
		7'd9: data <= {6'b100011, 5'b00000, 5'b01000, 16'b0000000000000100};
		7'd10: data <= {6'b000000, 5'b10001, 5'b10011, 5'b01001, 5'b00000, 6'b100000};
		7'd11: data <= {6'b000000, 5'b01000, 5'b10001, 5'b01010, 5'b00000, 6'b100000};
		7'd12: data <= {6'b100011, 5'b00000, 5'b01000, 16'b0000000000001000};
		7'd13: data <= {6'b000000, 5'b01000, 5'b10001, 5'b01010, 5'b00000, 6'b100000};
		7'd14: data <= {6'b100011, 5'b00000, 5'b01000, 16'b0000000000000100};
		7'd15: data <= {6'b101011, 5'b00000, 5'b01000, 16'b0000000000001100};
		7'd16: data <= {6'b000011, 26'b00000000000000000000010010};
		7'd17: data <= {6'b000100, 5'b10010, 5'b01000, 16'b0000000000000001};
		7'd18: data <= {6'b000000, 5'b11111, 5'b00000, 5'b00000, 5'b00000, 6'b001000};
		7'd19: data <= {6'b000010, 26'b00000000000000000000010011};
	   default:	data <= 32'h0000_0000;
	endcase
endmodule
