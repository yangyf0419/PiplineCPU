// rom_test3.v
//`timescale 1ns/1ps

module ROM_3 (addr,data);
    input [31:0] addr;
    output [31:0] data;
    reg [31:0] data;
    localparam ROM_SIZE = 32;
    reg [31:0] ROM_DATA[ROM_SIZE-1:0];

    always@(*)
        case(addr[9:2])   //Address Must Be Word Aligned.
            8'd0: data <= {6'b001000, 5'b00000, 5'b11111, 16'b0000000000000010};
            8'd1: data <= {6'b000000, 5'b11111, 5'b00000, 5'b00000, 5'b00000, 6'b001000};
            8'd2: data <= {6'b001111, 5'b00000, 5'b01000, 16'b0000000011111111};
            8'd3: data <= {6'b001000, 5'b01000, 5'b01001, 16'b0000000100000001};
            8'd4: data <= {6'b000000, 5'b00000, 5'b01001, 5'b10000, 5'b01000, 6'b000010};
            8'd5: data <= {6'b000000, 5'b00000, 5'b10000, 5'b10001, 5'b10000, 6'b000000};
            8'd6: data <= {6'b000000, 5'b00000, 5'b10001, 5'b10010, 5'b01100, 6'b000011};
            8'd7: data <= {6'b000000, 5'b10001, 5'b10010, 5'b10011, 5'b00000, 6'b101010};
            8'd8: data <= {6'b000000, 5'b10011, 5'b00000, 5'b10100, 5'b00000, 6'b100010};
            8'd9: data <= {6'b000110, 5'b10100, 5'b00000, 16'b0000000000000010};
            8'd10: data <= {6'b000000, 5'b10100, 5'b10011, 5'b10100, 5'b00000, 6'b100011};
            8'd11: data <= {6'b000011, 26'b00000000000000000000001001};
            8'd12: data <= {6'b000001, 5'b10100, 5'b00000, 16'b0000000000000011};
            8'd13: data <= {6'b001001, 5'b10100, 5'b10100, 16'b1111111111111111};
            8'd14: data <= {6'b000000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 6'b000000};
            8'd15: data <= {6'b000000, 5'b11111, 5'b00000, 5'b00000, 5'b00000, 6'b001000};
            8'd16: data <= {6'b000111, 5'b10100, 5'b00000, 16'b0000000000001001};
            8'd17: data <= {6'b000000, 5'b10100, 5'b01001, 5'b10100, 5'b00000, 6'b100001};
            8'd18: data <= {6'b000000, 5'b10100, 5'b10010, 5'b10100, 5'b00000, 6'b100110};
            8'd19: data <= {6'b000000, 5'b10100, 5'b10010, 5'b10100, 5'b00000, 6'b100111};
            8'd20: data <= {6'b001100, 5'b10100, 5'b10100, 16'b0000000100001111};
            8'd21: data <= {6'b001011, 5'b10010, 5'b01010, 16'b0000000000000011};
            8'd22: data <= {6'b001010, 5'b10010, 5'b01011, 16'b0000000000000010};
            8'd23: data <= {6'b000000, 5'b01011, 5'b10010, 5'b01011, 5'b00000, 6'b100101};
            8'd24: data <= {6'b000000, 5'b01011, 5'b10100, 5'b10100, 5'b00000, 6'b100100};
            8'd25: data <= {6'b000010, 26'b00000000000000000000010000};
            8'd26: data <= {6'b001000, 5'b00000, 5'b01100, 16'b0000000001011100};
            8'd27: data <= {6'b101011, 5'b01100, 5'b10010, 16'b0000000000000100};
            8'd28: data <= {6'b000100, 5'b10100, 5'b10100, 16'b0000000000000001};
            8'd29: data <= {6'b100011, 5'b01100, 5'b01101, 16'b0000000000000100};
            8'd30: data <= {6'b000101, 5'b10010, 5'b01101, 16'b1111111111111110};
            8'd31: data <= {6'b000000, 5'b01100, 5'b00000, 5'b11111, 5'b00000, 6'b001001};
            default: data <= 32'h80000000;
        endcase
endmodule


