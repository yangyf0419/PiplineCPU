// rom_test3.v
//`timescale 1ns/1ps

module ROM_3 (addr,data);
    input [31:0] addr;
    output [31:0] data;
    reg [31:0] data;
    localparam ROM_SIZE = 32;
    reg [31:0] ROM_DATA[ROM_SIZE-1:0];

    always@(*)
        case(addr[9:2])   //Address Must Be Word Aligned.
            // lui $t0, -256 # $t0 = 0x00ff0000
            8'd0:    data <= {6'b001111, 5'b00000, 5'b01000, 16'b1111111100000000};
            // addi $t1, $t0, 257 # $t1 = 0x00ff0101
            8'd1:    data <= {6'b001000, 5'b01000, 5'b01001, 16'b0000000100000001};
            // srl $s0, $t1, 8 # $s0 = 0x0000ff01
            8'd2:    data <= {6'b000000, 5'b00000, 5'b01001, 5'b10000, 5'b01000, 6'b000010};
            // sll $s1, $s0, 16 # $s1 = 0xff010000
            8'd3:    data <= {6'b000000, 5'b00000, 5'b10000, 5'b10001, 5'b10000, 6'b000000};
            // sra $s2, $s1, 12 # $s2 = 0xfffff010
            8'd4:    data <= {6'b000000, 5'b00000, 5'b10001, 5'b10010, 5'b01100, 6'b000011};
            // slt $s3, $s1, $s2 # $s3 = 0x00000001
            8'd5:    data <= {6'b000000, 5'b10001, 5'b10010, 5'b10011, 5'b00000, 6'b101010};
            // sub $s4, $s3, $zero # $s4 = 0x00000001
            8'd6:    data <= {6'b000000, 5'b10011, 5'b00000, 5'b10100, 5'b00000, 6'b100010};
            // L1:
            // blez $s4, L2
            8'd7:    data <= {6'b000110, 5'b10100, 5'b00000, 16'b0000000000000010};
            // subu $s4, $s4, $s3 # $s4 = 0
            8'd8:    data <= {6'b000000, 5'b10100, 5'b10011, 5'b10100, 5'b00000, 6'b100011}
            // jal L1
            8'd9:    data <= {6'b000011, 26'b00000000000000000000000111};
            // L2:
            // bltz $s4, L3
            8'd10:    data <= {6'b000001, 5'b10100, 5'b00000, 16'b0000000000000011}
            // addiu $s4, $s4, -1 # $s4 = -1
            8'd11:    data <= {6'b001001, 5'b10100, 5'b10100, 16'b1111111111111111}
            // nop
            8'd12:    data <= {6'b000000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 6'b000000}
            // jr $ra # j L2
            8'd13:    data <= {6'b000000, 5'b11111, 5'b00000, 5'b00000, 5'b00000, 6'b001000}
            // L3:
            // bgtz $s4, L4
            8'd14:    data <= {6'b000111, 5'b10100, 5'b00000, 16'b0000000000001001}
            // addu $s4, $s4, $t1 # $s4 = 0x00ff0100
            8'd15:    data <= {6'b000000, 5'b10100, 5'b01001, 5'b10100, 5'b00000, 6'b100001}
            // xor $s4, $s4, $s2 # $s4 = 0xff00f110
            8'd16:    data <= {6'b000000, 5'b10100, 5'b10010, 5'b10100, 5'b00000, 6'b100110}
            // nor $s4, $s4, $s2 # $s4 = 0x00000eef
            8'd17:    data <= {6'b000000, 5'b10100, 5'b10010, 5'b10100, 5'b00000, 6'b100111}
            // andi $s4, $s4, 271 # $s4 = 0x0000000f
            8'd18:    data <= {6'b001100, 5'b10100, 5'b10100, 16'b0000000100001111}
            // sltiu $t2, $s2, 3 # $t2 = 0x00000000
            8'd19:    data <= {6'b001011, 5'b10010, 5'b01010, 16'b0000000000000011}
            // slti $t3, $s2, 2 # $t3 = 0x00000001
            8'd20:    data <= {6'b001010, 5'b10010, 5'b01011, 16'b0000000000000010}
            // or $t3, $t3, $s2 # $t3 = 0xfffff011
            8'd21:    data <= {6'b000000, 5'b01011, 5'b10010, 5'b01011, 5'b00000, 6'b100101}
            // and $s4, $t3, $s4 # $s4 = 0x00000001
            8'd22:    data <= {6'b000000, 5'b01011, 5'b10100, 5'b10100, 5'b00000, 6'b100100}
            // j L3
            8'd23:    data <= {6'b000010, 26'b00000000000000000000001110}
            // L4:
            // addi $t4, $zero, 92 # $t4 = 0x0000005C
            8'd24:    data <= {6'b001000, 5'b00000, 5'b01100, 16'b0000000001011100}
            // sw $s2, 4($t4)
            8'd25:    data <= {6'b101011, 5'b01100, 5'b10010, 16'b0000000000000100}
            // beq $s4, $s4, L6
            8'd26:    data <= {6'b000100, 5'b10100, 5'b10100, 16'b0000000000000001}
            // lw $t5, 4($t4) # $t5 = 0xfffff010
            8'd27:    data <= {6'b100011, 5'b01100, 5'b01101, 16'b0000000000000100}
            // L6:
            // bne $s2, $t5, L5
            8'd28:    data <= {6'b000101, 5'b10010, 5'b01101, 16'b1111111111111110}
            // jalr $ra, $t4
            8'd29:    data <= {6'b000000, 5'b01100, 5'b00000, 5'b11111, 5'b00000, 6'b001001}
            default: data <= 32'h80000000;
        endcase
endmodule


